`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:10:01 05/16/2014 
// Design Name: 
// Module Name:    ColourControlLogic 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ColourControlLogic(
    input CLK,
	 input [1:0] MASTER_STATE,
    input [18:0] ADDR,
    input [7:0] CIN,
    output reg [7:0] COUT
    );


endmodule
